`ifndef _common_vh_
`define _common_vh_

// == supply rails ==
supply1 VCC;
supply0 GND;

`endif //_common_vh_
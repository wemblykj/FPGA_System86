`ifndef system86_system86_vh_
`define system86_system86_vh_

`include "common/common.vh"

`endif // system86_system86_vh_

entity system86 is
	generic
	(
	)
	port
	(
	
	);

end system86;

architecture rtl of system86 is

begin
end rtl;

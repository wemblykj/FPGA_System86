`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:       Paul Wightmore
// 
// Create Date:    11:16:41 05/12/2018 
// Design Name:    clut_subsystem
// Module Name:    system86/subsystem/videogen_subsystem.v 
// Project Name:   Namco System86 simulation
// Target Devices: 
// Tool versions: 
// Description:    videogen subsystem - 8-bit index to 4-bit RGB via CLUT
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
// License:        https://www.apache.org/licenses/LICENSE-2.0
//
//////////////////////////////////////////////////////////////////////////////////

module videogen_subsystem 
#(
)
(
    input CLK_6MD,
    input CLR,
    input [7:0] D,
    input BANK,
    output wire [3:0] RED,
    output wire [3:0] GREEN,
    output wire [3:0] BLUE,
    
    // == hardware abstraction - memory buses ==
    
    input wire [7:0] prom_3r_data,
    output wire [8:0] prom_3r_addr,
    output wire prom_3r_ce,
    
    input wire [3:0] prom_3s_data,
    output wire [8:0] prom_3s_addr,
    output wire prom_3s_ce
);
	
	assign BLUE = ls173_3v_d[7:4];
	assign GREEN = ls173_3u_d[7:4];
	assign RED = ls173_3t_d[7:4];
	
	wire [7:0] ls273_4u_d;
	ls273 ls273_4u(
		.CLK(CLK_6MD),
		.CLR(CLR),
		.D(D),
		.Q(ls273_4u_d)
		);
	
	wire [7:0] ls173_3v_d;
	ls173 ls173_3v(
		.CLK(CLK_6MD),
		.CLR(CLR),
		.D({prom_3s_data, 3'b0}),
		.Q(ls173_3v_d)
		);
		
	wire [7:0] ls173_3u_d;
	ls173 ls173_3u(
		.CLK(CLK_6MD),
		.CLR(CLR),
		.D({prom_3r_data[7:4], 3'b0}),
		.Q(ls173_3u_d)
		);
		
	wire [7:0] ls173_3t_d;
	ls173 ls173_3t(
		.CLK(CLK_6MD),
		.CLR(CLR),
		.D({prom_3r_data[3:0], 3'b0}),
		.Q(ls173_3t_d)
		);
		
	// == hardware abstraction - memory buses ==
    
	assign prom_3r_addr = {BANK, ls273_4u_d};
	assign prom_3r_ce = 1;
    
	assign prom_3s_addr = {BANK, ls273_4u_d};
	assign prom_3s_ce = 1;
    	
endmodule


`ifndef _rthunder_vh_
`define _rthunder_vh_
`include "roms.vh"

`define RTHUNDER "rthunder"

`define ROM_3R `MAKE_ROM_PATH(`RTHUNDER, "rtl-1.3r")
`define ROM_3S `MAKE_ROM_PATH(`RTHUNDER, "rt1-2.3s")


`define ROM_4R `MAKE_ROM_PATH(`RTHUNDER, "rt1_5.4r")
`define ROM_4S `MAKE_ROM_PATH(`RTHUNDER, "rt1_6.4s")
`define ROM_4V `MAKE_ROM_PATH(`RTHUNDER, "rt1-3.4v")

`define ROM_5V `MAKE_ROM_PATH(`RTHUNDER, "rt1-4.5v")

`define ROM_6U `MAKE_ROM_PATH(`RTHUNDER, "rt1-5.6u")

`define ROM_7R `MAKE_ROM_PATH(`RTHUNDER, "rt1_7.7r")
`define ROM_7S `MAKE_ROM_PATH(`RTHUNDER, "rt1_8.7s")

`define ROM_9C `MAKE_ROM_PATH(`RTHUNDER, "rt3_1b.9c")

`define ROM_12C `MAKE_ROM_PATH(`RTHUNDER, "rt3_2b.12c")
`define ROM_12D `MAKE_ROM_PATH(`RTHUNDER, "rt3_3.12d")



`endif //_rthunder_vh_
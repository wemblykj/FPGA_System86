`ifndef _rthunder_vh_
`define _rthunder_vh_
`include "roms.vh"

`define RTHUNDER "rthunder"

`define ROM_3R `MAKE_ROM_PATH(`RTHUNDER, "rtl-1.3r")
`define ROM_3S `MAKE_ROM_PATH(`RTHUNDER, "rt1-2.3s")

`endif //_rthunder_vh_
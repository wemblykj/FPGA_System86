`ifndef _common_vh_
`define _common_vh_

`define STRINGIFY(x) `"x`"

`endif //_common_vh_

library ieee;
use ieee.std_logic_1164.all;

entity system86 is

end system86;

architecture rtl of system86 is

begin
end rtl;

// This module is designed for 640x480 with a 25 MHz input clock.
`include "../../../../../../../lib/video_lib/rtl/VGA_Sync_Pulses.v"
`ifndef common_common_vh_
`define common_common_vh_

`define STRINGIFY(x) `"x`"

`endif // common_common_vh_


entity mc68a09e is
	generic
	(
	)
	port
	(
	
	);

end mc68a09e;

architecture rtl of mc68a09e is

begin
end rtl;
